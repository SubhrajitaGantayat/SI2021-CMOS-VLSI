***** Spice Netlist for Cell 'LAB9_inv' *****

************** Module LAB9_inv **************
m2 vout vin vdd vdd scmosp w='0.6u' l='0.4u' m='1' 
m1 vout vin gnd gnd scmosn w='0.6u' l='0.4u' m='1' 


.end

